module top
#(
  // Parameter list
 )
(
  // Port list
  /* Fill in inputs and outputs to module */
);

  counter
   #(
     .CYCLES_PER_COUNT ( 4 )
    )
  counter_i
    (
      /* Connect inputs and outputs of counter to
       * top module inputs and outputs */
    );

endmodule
